package fifo_pkg;
	`include "transaction.sv"
	`include "gen.sv"
	`include "drive.sv"
	`include "monitor.sv"
	`include "scoreboard.sv"
endpackage
