package fifo_pkg;
	`include "transaction.sv"
	`include "fifogenerator.sv"
	`include "fifodriver.sv"
	`include "fifomonitor.sv"
	`include "fifoscoreboard.sv"
endpackage
