/**********************************************************************/
/* ECE -593 FUNDAMENTALS OF PRESILICON VALIDATION                     */
/*				FINAL PROJECT										  */		
/* Authors : Achyuth Krishna Chepuri                                  */
/*			 Amrutha Regalla                                          */
/* 			 Sai Sri Harsha Atmakuri                                  */
/*			 Sathwik Reddy Madireddy                                  */ 
/**********************************************************************/

/*Driver module is responsible for converting transaction level stimuli generated by sequencer 
in signals and driving the actual interface. Build phase, connect phase and run phase are used to 
connect components and perform various actions.*/

class fifo_driver extends uvm_driver #(fifo_sequence_item);
`uvm_component_utils(fifo_driver)
virtual uvm_fifo vif;	
fifo_sequence_item item;

function new(string name ="fifo_driver",uvm_component parent);
		super.new (name,parent);
		`uvm_info("DRIVER CLASS", "fifo Driver",UVM_LOW)
endfunction
	
/******* BUILD PHASE *******/
function void build_phase (uvm_phase phase);
	super.build_phase(phase);
	`uvm_info("Driver Class", "Build Phase!",UVM_LOW)
	/*uvm_config_db is like central data base to store and retrieve various signals and interface*/
	if(!(uvm_config_db #(virtual uvm_fifo)::get(this,"*","vif",vif))) 
	begin
		`uvm_error("Driver Class", "Failed")
	end
endfunction


/******* CONNECT PHASE ******/
function void connect_phase(uvm_phase phase);
	super.connect_phase(phase);
	`uvm_info("Driver Class", "Connect Phase!",UVM_LOW)
endfunction

/******** RUN PHASE *******/
task run_phase(uvm_phase phase);
	super.run_phase(phase);
	`uvm_info("Driver Class", "Inside run Phase!",UVM_LOW)
	forever 
	 begin
		item = fifo_sequence_item#(8,9,512)::type_id::create("item");
		seq_item_port.get_next_item(item);
		drive(item);
		seq_item_port.item_done();
	 end
endtask

/******* DRIVE PHASE **********/
task drive(fifo_sequence_item item);
		begin
			if (!item.wrst & !item.rrst) begin
			vif.wrst <= item.wrst;
			vif.rrst <= item.rrst;
		end
		else begin
			if(item.winc & !item.rinc)
			  begin
			  vif.wrst <= item.wrst;
				vif.rrst <= item.rrst;
				vif.winc <= item.winc;
				vif.rinc <= item.rinc;
				vif.data_in <= item.data_in;
				@(posedge vif.wclk);			
				`uvm_info("DRIVER_WRITE",$sformatf("Burst Dtails:time=%0d,winc=%d,rinc=%d,data_in=%d,full=%0d,half_full=%0d,empty=%0d,half_empty=%0d,wr_addr=%d",$time,vif.winc,vif.rinc,vif.data_in,vif.full,vif.half_full,vif.empty,vif.half_empty,vif.wr_addr),UVM_LOW) 
				
			  end
			if(item.rinc & !item.winc)
			  begin
			    vif.wrst <= item.wrst;
				vif.rrst <= item.rrst;
				vif.rinc <= item.rinc;
				vif.winc <= item.winc;
				vif.data_in <= item.data_in;
				@(posedge vif.rclk);
				`uvm_info("DRIVER_READ",$sformatf("Burst Dtails:time=%0d,winc=%d,rinc=%d,data_out=%d,full=%0d,half_full=%0d,empty=%0d,half_empty=%0d,rd_addr=%d",$time,vif.winc,vif.rinc,vif.data_out,vif.full,vif.half_full,vif.empty,vif.half_empty,vif.rd_addr),UVM_LOW)
			    
			  end
			  
		end
	end
endtask

endclass