//Driver Code
